module fsm (
    input b_in,                 // 디바운싱된 버튼 입력
    input clk,                  // 시스템 클럭
    input rst_n,                // 리셋
    output reg [3:0] led_out    // 최종 LED 출력
);
    
    reg [1:0] state, next_state;
    parameter s0 = 2'b00, s1 = 2'b01, s2 = 2'b10, s3 = 2'b11;


    // --- 4. 엣지 검출 로직 (기존과 동일) ---
    reg b_in_prev;
    wire b_in_falling_edge;
    always @(posedge clk) begin
        b_in_prev <= b_in;
    end
    assign b_in_falling_edge = b_in_prev && !b_in;
    

    // --- 5. FSM 로직 수정 ---
    // 블록 1: 다음 상태 결정 (조합 회로)
    always @(*) begin
        next_state = state;
        // 버튼 하강 엣지가 감지될 때만 상태 변경
        if (b_in_falling_edge) begin
            case (state)
                s0: next_state = s1;
                s1: next_state = s2;
                s2: next_state = s3;
                s3: next_state = s0;
                default: next_state = s0;
            endcase
        end
    end

    // 블록 2: 상태 및 출력 업데이트 (순차 회로)
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= s0;
            led_out <= 4'b0001;
        end else begin
            state <= next_state;
            
            case (state)
                s0: led_out <= 4'b0001;
                s1: led_out <= 4'b0011;
                s2: led_out <= 4'b0111;
                s3: led_out <= 4'b1111;
                default: led_out <= 4'b0001;
            endcase
        end
    end

endmodule